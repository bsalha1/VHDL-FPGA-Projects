library ieee;
use ieee.std_logic_1164.all;

entity cpu is
end cpu;

architecture cpu_arch of cpu is
    signal address_bus : std_logic_vector(31 downto 0);
    
begin

end cpu_arch ;